// Code your design here

interface dut_if;

endinterface


module dut(dut_if dif);

endmodule
